module bin2bcd #(//????????
 parameter INPUT_WIDTH = 6,//??bit?????BCD??????????2^????-1
 parameter DECIMAL_DIGITS = 2//BCD??????????
 )(
 input i_Clock,//?????
 input [INPUT_WIDTH - 1 : 0] i_Binary,//??bit????
 input i_Start,//???????
 output [DECIMAL_DIGITS * 4 - 1 : 0] o_BCD,//???bit???????BCD????????????bit
 output o_DV//??????
 );


 parameter s_IDLE = 3'b000, s_SHIFT = 3'b001, s_CHECK_SHIFT_INDEX = 3'b010, s_ADD = 3'b011,//?????????????????
    s_CHECK_DIGIT_INDEX = 3'b100, s_BCD_DONE = 3'b101;

 reg [2:0] r_SM_Main = s_IDLE;//????????????????
   
  // The vector that contains the output BCD???????????????BCD??bit?
 reg [DECIMAL_DIGITS*4 - 1 : 0] r_BCD = 0;
    
  // The vector that contains the input binary value being shifted.?????????bit?
  reg [INPUT_WIDTH-1:0] r_Binary = 0;
      
  // Keeps track of which Decimal Digit we are indexing??????????BCD??
  reg [DECIMAL_DIGITS-1:0] r_Digit_Index = 0;
    
  // Keeps track of which loop iteration we are on.??????
  // Number of loops performed = INPUT_WIDTH???????????
  reg [7:0] r_Loop_Count = 0;
 
  wire [3:0] w_BCD_Digit;//??BCD???????
 reg r_DV = 1'b0;//?????????                      
    
  always @(posedge i_Clock) begin//?????????
      case (r_SM_Main)//?????????r_SM_Main??
  
        // Stay in this state until i_Start comes along????????????
        s_IDLE :
          begin
            r_DV <= 1'b0;
             
            if (i_Start == 1'b1)//?????????????bit?
              begin
                r_Binary  <= i_Binary;//r????????remain ?????
                r_SM_Main <= s_SHIFT;//???????
                r_BCD     <= 0;
              end
            else
              r_SM_Main <= s_IDLE;//???????????
          end
                 
  
        // Always shift the BCD Vector until we have shifted all bits through
        // Shift the most significant bit of r_Binary into r_BCD lowest bit.
        s_SHIFT :
          begin
            r_BCD     <= r_BCD << 1;
            r_BCD[0]  <= r_Binary[INPUT_WIDTH-1];//?binary????BCD?????
            r_Binary  <= r_Binary << 1;//binary??1Bit
            r_SM_Main <= s_CHECK_SHIFT_INDEX;//?????????
          end          
         
  
        // Check if we are done with shifting in r_Binary vector
        s_CHECK_SHIFT_INDEX :
          begin
            if (r_Loop_Count == INPUT_WIDTH-1)
              begin
                r_Loop_Count <= 0;//??????
                r_SM_Main    <= s_BCD_DONE;//????
              end
            else
              begin
                r_Loop_Count <= r_Loop_Count + 1;//??????
                r_SM_Main    <= s_ADD;//?????+3??
              end
          end
                 
  
        // Break down each BCD Digit individually.  Check them one-by-one to
        // see if they are greater than 4.  If they are, increment by 3.
        // Put the result back into r_BCD Vector.  
        s_ADD :
          begin
            if (w_BCD_Digit > 4)//??BCD???????????4
              begin                                     
                r_BCD[(r_Digit_Index*4)+:4] <= w_BCD_Digit + 3;//??4????????????3
              end
             
            r_SM_Main <= s_CHECK_DIGIT_INDEX; //?????BCD??????
          end       
         
         
        // Check if we are done incrementing all of the BCD Digits
        s_CHECK_DIGIT_INDEX :
          begin
            if (r_Digit_Index == DECIMAL_DIGITS-1)//??????
              begin
                r_Digit_Index <= 0;
                r_SM_Main     <= s_SHIFT;
              end
            else
              begin
                r_Digit_Index <= r_Digit_Index + 1;//BCD?????
                r_SM_Main     <= s_ADD;
              end
          end
         
  
  
        s_BCD_DONE :
          begin
            r_DV      <= 1'b1;//?????????????????????
            r_SM_Main <= s_IDLE;
          end
         
         
        default :
          r_SM_Main <= s_IDLE;//???????????
            
      endcase
    end // always @ (posedge i_Clock)  
 
   
  assign w_BCD_Digit = r_BCD[r_Digit_Index*4 +: 4];       
  assign o_BCD = r_BCD;                            

  assign o_DV  = r_DV;//??????????????????????????????
      			//????????????????????????????????
endmodule // Binary_to_BCD